`timescale 1 ps / 1 ps
// Instruction  Memory
module Inst_mem (
	Addr,
	clk,
	rst,
	q);

	input	[7:0]  Addr;
	input	  clk, rst;
	output	[15:0]  q;

	reg [7:0] ram [0:255]; //2 ^ 10 = 1024
	wire[15:0] addr_temp;
	always@(*)begin
		if(rst)begin
			ram[8'b00000000]=8'b00000000;
			ram[8'b00000001]=8'b00000000;
			ram[8'b00000010]=8'b00000000;
			ram[8'b00000011]=8'b00000000;
			ram[8'b00000100]=8'b01110000;
			ram[8'b00000101]=8'b00000000;
			ram[8'b00000110]=8'b11100000;
			ram[8'b00000111]=8'b11111111;
			ram[8'b00001000]=8'b11110000;
			ram[8'b00001001]=8'b00000111;
			ram[8'b00001010]=8'b11100000;
			ram[8'b00001011]=8'b00011111;
			ram[8'b00001100]=8'b11110000;
			ram[8'b00001101]=8'b11111111;
			ram[8'b00001110]=8'b11110100;
			ram[8'b00001111]=8'b11111111;
			ram[8'b00010000]=8'b01010000;
			ram[8'b00010001]=8'b00000000;
			ram[8'b00010010]=8'b01000100;
			ram[8'b00010011]=8'b00000000;
			ram[8'b00010100]=8'b10001100;
			ram[8'b00010101]=8'b00000000;
			ram[8'b00010110]=8'b11010000;
			ram[8'b00010111]=8'b11111111;
			ram[8'b00011000]=8'b01010000;
			ram[8'b00011001]=8'b00000000;
			ram[8'b00011010]=8'b11100000;
			ram[8'b00011011]=8'b11111111;
			ram[8'b00011100]=8'b10000011;
			ram[8'b00011101]=8'b00000000;
			ram[8'b00011110]=8'b10100000;
			ram[8'b00011111]=8'b00100100;
			ram[8'b00100000]=8'b00010001;
			ram[8'b00100001]=8'b00000000;
			ram[8'b00100010]=8'b10010000;
			ram[8'b00100011]=8'b00100110;
			ram[8'b00100100]=8'b00110001;
			ram[8'b00100101]=8'b00000000;
			ram[8'b00100110]=8'b01100000;
			ram[8'b00100111]=8'b00000000;
			ram[8'b00101000]=8'b10110000;
			ram[8'b00101001]=8'b00110100;
			ram[8'b00101010]=8'b10000011;
			ram[8'b00101011]=8'b00000000;
			ram[8'b00101100]=8'b10100100;
			ram[8'b00101101]=8'b00110000;
			ram[8'b00101110]=8'b10010000;
			ram[8'b00101111]=8'b00010000;
			ram[8'b00110000]=8'b10010000;
			ram[8'b00110001]=8'b00000100;
			ram[8'b00110010]=8'b00000000;
			ram[8'b00110011]=8'b00000000;
			ram[8'b00110100]=8'b11010000;
			ram[8'b00110101]=8'b00011111;
			ram[8'b00110110]=8'b10001001;
			ram[8'b00110111]=8'b00000000;
			ram[8'b00111000]=8'b11110100;
			ram[8'b00111001]=8'b00000001;
			ram[8'b00111010]=8'b00100001;
			ram[8'b00111011]=8'b00000000;
			ram[8'b00111100]=8'b11100000;
			ram[8'b00111101]=8'b00011111;
			ram[8'b00111110]=8'b10000110;
			ram[8'b00111111]=8'b00000000;
			ram[8'b01000000]=8'b11000000;
			ram[8'b01000001]=8'b00000000;
		end
	end
	assign addr_temp = (Addr>>1)<<1;
	assign q = {ram[addr_temp+1],ram[addr_temp]};
endmodule
